package pkg;
  import uvm_pkg::*;
  `include "sequence_item.sv"
  `include "sequence.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include "test.sv"
  
  // Add other files as you create them
endpackage